module signed_adder
(
	input signed [3:0] a,
	input 		 [3:0] b,
	input			   cin,
	output signed [5:0] sum
);

	assign sum = {a[3], a} < {1'b0, b};
endmodule
